My Test Circuit
* Generated netlist

VW1 0 nodeA SIN(0 5 1k 0 0 0)
R1 nodeA nodeB 1k
R2 nodeB 0 1k

* Labeled Nodes:
* Node 0 = 0
* Node 2 = nodeA
* Node 3 = nodeB

* Simulation Options
.option TEMP=27
.option TNOM=27

* Analysis Command
.op

* Control block for batch execution
.control
set wr_vecnames  * Ensure header is printed for table
run
print v(nodeA) v(nodeB)
wrdata transient_data.txt v(nodeA) v(nodeB)
.endc

.end