MOSFET Switched Resistor

*the purpose of this circuit is to gain familiarity with MOSFETS and using dummy voltage sources to measure current. All values were selected semi-arbitrarily.

VCC 1 0 DC 12
R1 1 2 10

Vmeas 2 3
*Vmeas is a 0v source i.e. short. This acts like an ideal ammeter allowing current to be measured.

M1 3 4 0 0 MMOD
*MOSFET M1 has drain connected to node 3, gate connected to node 4, source grounded, and substrate grounded. Note: source and substrate are almost always connected to the same node.

Vpwm 4 0 pulse(0 10 0 1ns 1ns 2ms 4ms)
*Vpwm is a pulse train with 0 offset, pulsed value of 10v, 0 time delay, 1ns rise time, 1ns fall time, 2ms pulse width, and 4ms period.

.tran 1ns 10ms

.model MMOD NMOS
*defines model MMOD as an N-channel MOSFET with default parameters

.control
run

plot i(Vmeas)
*plots the currect through Vmeas (our pseudo ammeter)

.endc
.end
