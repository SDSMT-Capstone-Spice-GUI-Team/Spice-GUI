MOSFET Switched Motor

*the purpose of this circuit was to represent a motor with current controlled by a MOSFET driven by a pulse-width modulation (pwm) signal. motor is represented by 1000ohm resistance and 5H inductance with back EMF being ignored. all values were chosen semi-arbitrarily.

VCC 1 0 DC 12

R1 1 2 1000
*R1 represents motor resistance

L1 2 3 5
*inductor L1 is connected to nodes 2 and 3 with 5H inductance. L1 represents motor inductance

Vmeas 3 4
*Vmeas is used as an ammeter to measure current through the motor

D1 4 1 DMOD
M1 4 5 0 0 MMOD
Vpwm 5 0 pulse(0 10 0 1ns 1ns 1ms 2ms)

.tran 1ns 10ms
.model DMOD D
.model MMOD NMOS
.control
run
plot i(Vmeas)
.endc
.end
